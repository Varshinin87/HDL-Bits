// Description: This is a simple pass-through module where the input signal is directly assigned to the output.

module top_module( input in, output out );  

    // Assign the input 'in' directly to the output 'out'
    assign out = in;  

endmodule  
