module top_module (
    input in,    // Single-bit input
    output out   // Single-bit output
);

assign out = in;  // Assign the input directly to the output

endmodule
