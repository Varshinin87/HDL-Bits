module top_module (
    output out   // Single-bit output
);

assign out = 1'b0;  // Assign a constant 0 to the output

endmodule
