module top_module( input in, output out );  

    // Assign the input 'in' directly to the output 'out'
    assign out = in;  

endmodule  
