module top_module (
    input a,        // 1-bit input 'a' to the top module
    input b,        // 1-bit input 'b' to the top module
    output out      // 1-bit output 'out' from the top module
);

    // Instantiate the submodule 'mod_a' named 'instance1'
    // Connect inputs 'a' and 'b' from the top module to 'mod_a' instance
    // The output of 'mod_a' is connected to 'out' in the top module
    mod_a instance1 (
        .in1(a),        // Connect 'a' input to 'a' input of mod_a
        .in2(b),        // Connect 'b' input to 'b' input of mod_a
        .out(out)     // Connect 'out' output of mod_a to the 'out' of the top module
    );            

endmodule
